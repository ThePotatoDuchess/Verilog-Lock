module LCDdisp (clk,num,Lclk,Lrst,Ldata,Lms,Lss);
input clk;
input [2:0]num;
output Lclk,Lrst,Ldata,Lms,Lss;
parameter SIZE = 8192;
wire [0:SIZE] img;
reg [14:0] pos;
reg Ldata;
reg Lclk;
reg Lrst;
reg store;

initial
begin
store = 1;
end


imgDAT i1 (store,img);

always @(posedge clk)
begin
		if(pos<SIZE &~Lrst)
		begin
			Ldata = img[pos];
			Lclk = ~Lclk;
			pos = pos+1;
		end
		else if (~(store==num))
		begin
			pos = 0;
			Lrst = 1;
			store = num;
		end
		else if (Lrst)
		begin
		Lrst = 0;
		
		end

end


endmodule


module imgDAT(num,img);
input [2:0] num;
output [0:8192] img;
reg img;

always @(num)
begin
	case(num)
	2'b01 : img = 8192'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000100010001000100010001000100010001000100010001000000000001000100010001000100010001000100010001000100000000000000010001000100000000000000000000000100010001000000000000000100010001000100010001000100010001000100010000000000000001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000001000100010001000100010001000100010001000100010000000000010001000100010001000100010001000100010001000000000000000100010001000000000000000000010001000100010000000000000001000100010001000100010001000100010001000100000000000000010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000010001000100010001000100010001000100010001000100000000000100010001000100010001000100010001000100010000000000000001000100010000000000000001000100010001000100000000000000010001000100010001000100010001000100010001000000000000000100010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000100010001000000000000000000000000000100010001000000000001000100010000000000000000000000000000000000000000000000010001000100000000000100010001000100010000000000000000000100010001000000000000000000000000000000000000000000000001000100010000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000001000100010000000000000000000000000001000100010000000000010001000100000000000000000000000000000000000000000000000100010001000000010001000100010001000000000000000000000001000100010000000000000000000000000000000000000000000000010001000100000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000010001000100000000000000000000000000010001000100000000000100010001000000000000000000000000000000000000000000000001000100010001000100010001000100000000000000000000000000010001000100000000000000000000000000000000000000000000000100010001000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000100010001000000000000000000000000000100010001000000000001000100010000000000000000000000000000000000000000000000010001000100010001000100010000000000000000000000000000000100010001000100010001000100010001000100010000000000000001000100010000000000000000000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000001000100010000000000000000000000000001000100010000000000010001000100000000000000000000000000000000000000000000000100010001000100010001000000000000000000000000000000000001000100010001000100010001000100010001000100000000000000010001000100000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000010001000100000000000000000000000000010001000100000000000100010001000000000000000000000000000000000000000000000001000100010001000100010000000000000000000000000000000000010001000100010001000100010001000100010001000000000000000100010001000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000100010001000000000000000000000000000100010001000000000001000100010000000000000000000000000000000000000000000000010001000100010001000100010000000000000000000000000000000100010001000000000000000000000000000000000000000000000001000100010000000000000000000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000001000100010000000000000000000000000001000100010000000000010001000100000000000000000000000000000000000000000000000100010001000100010001000100010000000000000000000000000001000100010000000000000000000000000000000000000000000000010001000100000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000010001000100000000000000000000000000010001000100000000000100010001000000000000000000000000000000000000000000000001000100010000000100010001000100010000000000000000000000010001000100000000000000000000000000000000000000000000000100010001000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000100010001000000000000000000000000000100010001000000000001000100010000000000000000000000000000000000000000000000010001000100000000000100010001000100010000000000000000000100010001000000000000000000000000000000000000000000000001000100010000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100010001000100010001000100010001000000000001000100010001000100010001000100010001000100010000000000010001000100010001000100010001000100010001000000000000000100010001000000000000000100010001000100010000000000000001000100010001000100010001000100010001000100000000000000010001000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000100010001000100010001000100010000000000010001000100010001000100010001000100010001000100000000000100010001000100010001000100010001000100010000000000000001000100010000000000000000000100010001000100000000000000010001000100010001000100010001000100010001000000000000000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010001000100010001000100010001000100000000000100010001000100010001000100010001000100010001000000000001000100010001000100010001000100010001000100000000000000010001000100000000000000000000000100010001000000000000000100010001000100010001000100010001000100010000000000000001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000000000100010001000100010001000100010001000100010001000000000001000100010001000100010001000100010001000000000000000000010001000100010001000100010001000100010001000100000000000100010001000100010001000100010001000100010000000000000001000100010001000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000001000100010001000100010001000100010001000100010000000000010001000100010001000100010001000100010001000000000000000100010001000100010001000100010001000100010001000000000001000100010001000100010001000100010001000100000000000000010001000100010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000010001000100010001000100010001000100010001000100000000000100010001000000000000000000000000000100010001000000000001000100010001000100010001000100010001000100010000000000010001000100010001000100010001000100010001000000000000000100010001000100010001000100010001000100010001000000000000000000010001000100010000000000000000000000000000000100010001000100010000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000001000100010000000000000000000000000000000100010000000000000000000000000001000100010001000000000000000000000000000100010001000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000010001000100010001000100000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000010001000100000000000000000000000000000001000100000000000000000000000000010001000100010000000000000000000000000001000100010000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000000001000100010001000000000000000000000001000100010001000100010001000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000100010001000000000000000000000000000000010001000000000000000000000000000100010001000100000000000000000000000000010001000100000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000010001000100010000000000000000000100010001000100010001000100010000000000000000000000000000000000000000000100010001000100010001000100010001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000001000100010000000000000000000000000000000100010000000000000000000000000001000100010001000000000000000000000000000100010001000100010001000100010001000100000000000000000001000100010001000100010001000100010001000100010000000000000000000000000000000000000000000000000001000100010001000000010001000100000000000000000000000000000000000000000001000100010001000100010001000100010001000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000010001000100000000000000000000000000010001000100000000000000000000000000010001000100010000000000000000000000000001000100010001000100010001000100010001000000000000000000010001000100010001000100010001000100010001000100000000000000000000000000000000000000000000000000010001000100000000000100010001000000000000000000000000000000000000000000010001000100010001000100010001000100010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000100010001000100010001000100010001000100010000000000000000000000000000000100010001000100000000000000000000000000010001000100010001000100010001000100010000000000000000000100010001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000100010001000100010001000100010001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000001000100010001000100010001000100010001000000000000000000000000000000000001000100010001000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000000000000000000000000000001000100010001000100010001000100000000000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000010001000100000000000100010001000000000000000000000000000000000000000000010001000100010000000000000000000000000001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000000000001000100010001000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000010001000100010001000100010000000100010000000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000100010001000000000000000100010001000000000000000000000000000000000000000100010001000100000000000000000000000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000010001000100010000000000000000000000000000000000000001000100010000000000000000000000000000000000000000000100010001000100010001000100000001000100000001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000001000100010000000000000000000100010001000000000000000000000000000000000001000100010001000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000000000000100010001000100000000000000000000000000000000000000010001000100000000000000000000000000000000000000000001000100010001000100010001000100000000000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000010001000100000000000000000000000100010001000000000000000100010001000100010001000100010001000100010001000000000001000100010001000100010001000100010001000100000000000000010001000100010001000100010001000100010001000100000000000000000001000100010001000000000000000000010001000100010001000100010001000100010001000100000000000000000000000000010001000100010001000100010001000000000001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000100010001000000000000000000000000000100010001000000000001000100010001000100010001000100010001000100010000000000010001000100010001000100010001000100010001000000000000000100010001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000100010001000100010001000100010001000100010001000000000000000000000000000100010001000100010001000100000000000000000001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000001000100010000000000000000000000000000000100010000000000010001000100010001000100010001000100010001000100000000000100010001000100010001000100010001000100010000000000000001000100010001000100010001000100010001000100010000000000000000000000000000000000000000000000000001000100010001000100010001000100010001000100010000000000000000000000000001000100010001000100010001000000000000000000010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010001000100000000000000000000000000010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100010001000000000000000000000000000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000100010001000100010001000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010001000100010001000100010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100010001000100010001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000100010001000100010001000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	endcase

end

endmodule